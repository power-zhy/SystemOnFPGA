`include "define.vh"


/**
 * UART RX part for receiving data only.
 * Author: Zhao, Hongyu  <power_zhy@foxmail.com>
 */
module uart_core_rx (
	input wire clk,  // main clock
	input wire rst,  // synchronous reset
	input wire [BAUD_DIV_WIDTH-1:0] baud_div,  // baud rate division, should be 10M/8/baudrate-1
	input wire [1:0] data_type,  // type for number of data bits, 00 for eight, 01 for seven, 10 for six, 11 for five
	input wire [1:0] stop_type,  // type for number of stop bits, 00 for one, 01 for one and a half, 10 for two
	input wire check_en,  // whether to use data checking or not
	input wire [1:0] check_type,  // data checking type, 00 for odd, 01 for even, 10 for mark, 11 for space
	input wire en,  // enable signal
	output reg [DATA_BITS_MAX-1:0] data,  // data received in
	output reg busy,  // busy flag
	output reg ack,  // data received acknowledge
	output reg err,  // data checking error
	// UART TX interface
	input wire rx
	);
	
	`include "function.vh"
	parameter
		CLK_FREQ = 100,  // main clock frequency in MHz, should be multiple of 10M
		BAUD_DIV_WIDTH = 8;  // width for baud rate division
	localparam
		DATA_BITS_MAX = 8,  // maximum data length for transmit
		STOP_BITS_MAX = 2,  // maximum stop flag length
		SAMPLE_COUNT = 8,
		SAMPLE_COUNT_WIDTH = GET_WIDTH(SAMPLE_COUNT-1),
		CLK_DIV = CLK_FREQ / 10,
		CLK_DIV_WIDTH = GET_WIDTH(CLK_DIV-1),
		TRANS_BITS_MAX = DATA_BITS_MAX + STOP_BITS_MAX,  // no need to store the start bit and last stop bit in current implement
		TRANS_BITS_WIDTH = GET_WIDTH(TRANS_BITS_MAX);
	
	reg check_bit;
	reg [TRANS_BITS_WIDTH-1:0] trans_bits;
	reg [TRANS_BITS_MAX-1:0] data_buf;
	reg [CLK_DIV_WIDTH-1:0] clk_count = 0;
	reg [BAUD_DIV_WIDTH-1:0] hns_count = 0;
	reg [SAMPLE_COUNT_WIDTH-1:0] sample_count = 0;
	reg [SAMPLE_COUNT_WIDTH-1:0] pos_count = 0;
	reg [SAMPLE_COUNT_WIDTH-1:0] neg_count = 0;
	reg [TRANS_BITS_WIDTH-1:0] bit_count = 0;
	
	always @(*) begin
		case (data_type)  // regard one and a half stop bits as one
			2'b00: case (stop_type)
				2'b10: trans_bits = check_en ? 4'd11 : 4'd10;
				default: trans_bits = check_en ? 4'd10 : 4'd9;
			endcase
			2'b01: case (stop_type)
				2'b10: trans_bits = check_en ? 4'd10 : 4'd9;
				default: trans_bits = check_en ? 4'd9 : 4'd8;
			endcase
			2'b10: case (stop_type)
				2'b10: trans_bits = check_en ? 4'd9 : 4'd8;
				default: trans_bits = check_en ? 4'd8 : 4'd7;
			endcase
			2'b11: case (stop_type)
				2'b10: trans_bits = check_en ? 4'd8 : 4'd7;
				default: trans_bits = check_en ? 4'd7 : 4'd6;
			endcase
		endcase
	end
	
	always @(*) begin
		if (check_en) begin
			case (check_type)
				2'b00: begin
					case (data_type)
						2'b00: check_bit = ~(^data[7:0]);
						2'b01: check_bit = ~(^data[6:0]);
						2'b10: check_bit = ~(^data[5:0]);
						2'b11: check_bit = ~(^data[4:0]);
					endcase
				end
				2'b01: begin
					case (data_type)
						2'b00: check_bit = (^data[7:0]);
						2'b01: check_bit = (^data[6:0]);
						2'b10: check_bit = (^data[5:0]);
						2'b11: check_bit = (^data[4:0]);
					endcase
				end
				2'b10: check_bit = 1;
				2'b11: check_bit = 0;
			endcase
		end
		else begin
			check_bit = 0;
		end
	end
	
	reg checked;
	always @(*) begin
		case ({check_en, data_type})  // last stop bit is not in data_buf
			3'b000: case (stop_type)
				2'b10: {checked, data[7:0]} = {1'b0, data_buf[TRANS_BITS_MAX-2:TRANS_BITS_MAX-9]};
				default: {checked, data[7:0]} = {1'b0, data_buf[TRANS_BITS_MAX-1:TRANS_BITS_MAX-8]};
			endcase
			3'b001: case (stop_type)
				2'b10: {checked, data[7:0]} = {2'b0, data_buf[TRANS_BITS_MAX-2:TRANS_BITS_MAX-8]};
				default: {checked, data[7:0]} = {2'b0, data_buf[TRANS_BITS_MAX-1:TRANS_BITS_MAX-7]};
			endcase
			3'b010: case (stop_type)
				2'b10: {checked, data[7:0]} = {3'b0, data_buf[TRANS_BITS_MAX-2:TRANS_BITS_MAX-7]};
				default: {checked, data[7:0]} = {3'b0, data_buf[TRANS_BITS_MAX-1:TRANS_BITS_MAX-6]};
			endcase
			3'b011: case (stop_type)
				2'b10: {checked, data[7:0]} = {4'b0, data_buf[TRANS_BITS_MAX-2:TRANS_BITS_MAX-6]};
				default: {checked, data[7:0]} = {4'b0, data_buf[TRANS_BITS_MAX-1:TRANS_BITS_MAX-5]};
			endcase
			3'b100: case (stop_type)
				2'b10: {checked, data[7:0]} = {data_buf[TRANS_BITS_MAX-2:TRANS_BITS_MAX-10]};
				default: {checked, data[7:0]} = {data_buf[TRANS_BITS_MAX-1:TRANS_BITS_MAX-9]};
			endcase
			3'b101: case (stop_type)
				2'b10: {checked, data[7:0]} = {data_buf[TRANS_BITS_MAX-2], 1'b0, data_buf[TRANS_BITS_MAX-3:TRANS_BITS_MAX-9]};
				default: {checked, data[7:0]} = {data_buf[TRANS_BITS_MAX-1], 1'b0, data_buf[TRANS_BITS_MAX-2:TRANS_BITS_MAX-8]};
			endcase
			3'b110: case (stop_type)
				2'b10: {checked, data[7:0]} = {data_buf[TRANS_BITS_MAX-2], 2'b0, data_buf[TRANS_BITS_MAX-3:TRANS_BITS_MAX-8]};
				default: {checked, data[7:0]} = {data_buf[TRANS_BITS_MAX-1], 2'b0, data_buf[TRANS_BITS_MAX-2:TRANS_BITS_MAX-7]};
			endcase
			3'b111: case (stop_type)
				2'b10: {checked, data[7:0]} = {data_buf[TRANS_BITS_MAX-2], 3'b0, data_buf[TRANS_BITS_MAX-3:TRANS_BITS_MAX-7]};
				default: {checked, data[7:0]} = {data_buf[TRANS_BITS_MAX-1], 3'b0, data_buf[TRANS_BITS_MAX-2:TRANS_BITS_MAX-6]};
			endcase
		endcase
	end
	
	always @(posedge clk) begin
		ack <= 0;
		err <= 0;
		if (rst) begin
			clk_count <= 0;
			hns_count <= 0;
			sample_count <= 0;
			pos_count <= 0;
			neg_count <= 0;
			bit_count <= 0;
			data_buf <= 0;
		end
		else if (busy) begin
			if (clk_count != CLK_DIV-1) begin
				clk_count <= clk_count + 1'h1;
			end
			else begin
				clk_count <= 0;
				if (hns_count != baud_div) begin
					hns_count <= hns_count + 1'h1;
				end
				else begin
					hns_count <= 0;
					if (sample_count != SAMPLE_COUNT-1) begin
						if (rx)
							pos_count <= pos_count + 1'h1;
						else
							neg_count <= neg_count + 1'h1;
						sample_count <= sample_count + 1'h1;
					end
					else begin
						sample_count <= 0;
						pos_count <= 0;
						neg_count <= 0;
						/*if (bit_count != trans_bits) begin
							bit_count <= bit_count + 1'h1;
							data_buf <= {(pos_count > neg_count), data_buf[TRANS_BITS_MAX-1:1]};  // would not save the last stop bit
						end
						else begin
							bit_count <= 0;
							if (pos_count > neg_count && checked == check_bit)
								ack <= 1;
							else
								err <= 1;
						end*/
						if (bit_count == trans_bits-1'h1) begin
							ack <= 1;
							bit_count <= 0;
						end
						else begin
							bit_count <= bit_count + 1'h1;
						end
						data_buf <= {(pos_count > neg_count), data_buf[TRANS_BITS_MAX-1:1]};  // would not save the last stop bit
					end
				end
			end
		end
		else begin
			clk_count <= 0;
			hns_count <= 0;
			sample_count <= 0;
			pos_count <= 0;
			neg_count <= 0;
			bit_count <= 0;
			data_buf <= 0;
		end
	end
	
	reg rx_prev;
	always @(posedge clk) begin
		if (rst)
			rx_prev <= 0;
		else
			rx_prev <= rx;
	end
	
	localparam
		S_IDLE = 0,  // idle
		S_START = 1,  // receive and check start bit
		S_TRANS = 2;  // receive data
	
	reg [1:0] state = 0;
	reg [1:0] next_state;
	
	always @(*) begin
		next_state = S_IDLE;
		case (state)
			S_IDLE: begin
				if (en && rx_prev && ~rx)
					next_state = S_START;
				else
					next_state = S_IDLE;
			end
			S_START: begin
				if (bit_count == 1)
					if (data_buf[TRANS_BITS_MAX-1])  // invalid start bit
						next_state = S_IDLE;
					else
						next_state = S_TRANS;
				else
					next_state = S_START;
			end
			S_TRANS: begin
				if (ack || err)
					next_state = S_IDLE;
				else
					next_state = S_TRANS;
			end
		endcase
	end
	
	always @(posedge clk) begin
		if (rst)
			state <= 0;
		else
			state <= next_state;
	end
	
	always @(posedge clk) begin
		if (rst) begin
			busy <= 0;
		end
		else case (next_state)
			S_IDLE: begin
				busy <= 0;
			end
			default: begin
				busy <= 1;
			end
		endcase
	end
	
endmodule
