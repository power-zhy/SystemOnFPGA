// Memory Access Type
localparam
	MEM_TYPE_WORD  = 2'h0,
	MEM_TYPE_HALF  = 2'h1,
	MEM_TYPE_BYTE  = 2'h2;
